module two_input_and (
  input A,
  input B,
  output Y
);

  assign Y = A & B;

endmodule