module two_input_or (
  input A,
  input B,
  output Y
);

  assign Y = A | B;

endmodule