module two_input_xor (
  input A,
  input B,
  output Y
);

  assign Y = A ^ B;

endmodule